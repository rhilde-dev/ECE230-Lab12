module ripple_counter();




endmodule;